library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller is
	port (
		clk   : in std_logic;
		reset : in std_logic;
	);
end controller;

architecture controllerArch of controller is
begin

end controllerArch;
